module SlowClock(
	input wire clk, reset, 
	output reg clk_1Hz
);

reg [27:0] counter;

always@(posedge reset or posedge clk)
begin
    if (reset == 1'b1)
        begin
            clk_1Hz <= 0;
            counter <= 0;
        end
    else
        begin
            counter <= counter + 1;
            if ( counter == 4_000)
                begin
                    counter <= 0;
                    clk_1Hz <= clk_1Hz + 1;
                end
        end
end
endmodule   